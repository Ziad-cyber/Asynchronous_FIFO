module FIFO (
    
);
    
endmodule